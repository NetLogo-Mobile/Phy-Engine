module alu16_mov(
    input  wire [15:0] b,
    output wire [15:0] y
);
    assign y = b;
endmodule
